module main

import user_interface as ui	// Import our custom UI.

fn main()
{
    mut app := ui.App{}		//
    app.start()				// Create app instance and start it
}